--/*
--**********************************************************
--  Design Automation Course Homework (Spring, 2020 Semester)
--  Amirkabir University of Technology (Tehran Polytechnic)
--  Department of Computer Engineering (CE-AUT)
--  https://ce.aut.ac.ir
--  Created by TA (ali[dot]mohammadpour[at]ac[dot]ir)
--  *******************************************************
--  Student ID  : XXXXXXX
--  Student Name: -----------------
--  Student Mail: -----------------
--  *******************************************************
--  Module: ProblemSet 4, Problem 4, Squence Detector 
--  *******************************************************
--  Additional Comments:
--*/

library ieee;
use ieee.std_logic_1164.all;

entity sequence_detector is
	port (
		clock    : in  std_logic ;
		reset    : in  std_logic ;
		din      : in  std_logic ;
		detected : out std_logic ) ;
end sequence_detector;

architecture sequence_detector_arch of sequence_detector is

	-- write your code, module is a fsm (johnson)

begin

	-- write your code here

end sequence_detector_arch;
