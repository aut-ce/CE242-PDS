--/*
--**********************************************************
--  Design Automation Course Homework (Spring, 2020 Semester)
--  Amirkabir University of Technology (Tehran Polytechnic)
--  Department of Computer Engineering (CE-AUT)
--  https://ce.aut.ac.ir
--  Designed TA (ali[dot]mohammadpour[at]ac[dot]ir)
--  *******************************************************
--  Student ID  : XXXXXXX
--  Student Name: -----------------
--  Student Mail: -----------------
--  *******************************************************
--  Module: ProblemSet 3, Problem 2, Section A
--  *******************************************************
--  Additional Comments:
--*/

library ieee;
use ieee.std_logic_1164.all;

entity piso is
	port (
		clk : in std_logic ;
		para_in : in std_logic_vector ;
		reset : in std_logic ;
		load : in std_logic ; 
		shift_en : in std_logic ; 
		ser_out : out std_logic) ;
end piso;

architecture piso_arc of piso is

begin

     -- write your code here

end  piso_arc;

