package riscv_types_pkg is
	
end package riscv_types_pkg;

package body riscv_types_pkg is

end package body riscv_types_pkg;


entity test is
end entity ;

architecture arch of test is

	-- use defined record type


begin

end architecture ;
