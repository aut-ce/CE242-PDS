--/*
--**********************************************************
--  Design Automation Course Homework (Spring, 2020 Semester)
--  Amirkabir University of Technology (Tehran Polytechnic)
--  Department of Computer Engineering (CE-AUT)
--  https://ce.aut.ac.ir
--  Designed TA (ali[dot]mohammadpour[at]ac[dot]ir)
--  *******************************************************
--  Student ID  : XXXXXXX
--  Student Name: -----------------
--  Student Mail: -----------------
--  *******************************************************
--  Module: ProblemSet 3, Problem 5
--  *******************************************************
--  Additional Comments:
--*/

library ieee;
use ieee.std_logic_1164.all;

entity problem_3_5 is
	port (
		time_x  : in aut_time_t ;
		time_y 	 : in aut_time_t ;
		operation	 : in std_logic ;
		time_o 	 : out aut_time_t );
end problem_3_5;

architecture problem_3_5_arc of problem_3 is

     -- write your code here

begin

     -- write your code here

end  problem_3_5_arc;

------------------------------------------------------
------------------------------------------------------

-- create new package and add time type to it.
-- in problem_3_5_arc use time type + and - opetations

