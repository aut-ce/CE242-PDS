library ieee;
use ieee.std_logic_1164.all;

library xil_defaultlib;
use xil_defaultlib.xpoint_pkg.all;

entity tanh is
	port (
		x    : in  xfixed(2 downto -3);
		outp : out std_logic_vector(15 downto 0));
end tanh;

architecture arc_lutx of tanh is
	type lookups is array (0 to 63) of std_logic_vector(15 downto 0);
	constant tanh_lookups : lookups := (
			"0011110000000000", "0011110000000000", "0011110000000000", "0011110000000000",
			"0011110000000000", "0011110000000000", "1011011010000000", "1011011010000000",
			"1011101000000000", "1011101000000000", "1011011000000000", "1011101000000000",
			"1011101000000000", "1011101000000000", "1011110000000000", "1011110000000000",
			"1011110000000000", "1011110000000000", "1011110000000000", "1011110000000000",
			"1011110000000000", "1011110000000000", "1011011010000000", "1011011010000000",
			"1011011010000000", "1011011010000000", "1011011010000000", "1011011010000000",
			"1011011010000000", "1011101000000000", "1011101000000000", "1011011000000000",
			"1011101000000000", "1011101000000000", "1011101000000000", "1011110000000000",
			"1011110000000000", "1011110000000000", "1011110000000000", "1011110000000000",
			"1011110000000000", "1011110000000000", "1011110000000000", "1011011010000000",
			"1011011010000000", "1011011010000000", "1011011010000000", "1011011010000000",
			"1011011010000000", "1011011010000000", "1011101000000000", "1011101000000000",
			"1011011000000000", "1011101000000000", "1011101000000000", "1011101000000000",
			"1011110000000000", "1011110000000000", "1011110000000000", "1011110000000000",
			"1011110000000000", "1011110000000000", "1011110000000000", "1011110000000000");

begin

	outp <= tanh_lookups(to_integer(unsigned(x)));

end arc_lutx;

architecture arc_hard of tanh is
	constant tanh_lookups : lookups := (
			"0011110000000000", "0011110000000000", "0011110000000000", "0011110000000000",
			"0011110000000000", "0011110000000000", "1011011010000000", "1011011010000000",
			"1011101000000000", "1011101000000000", "1011011000000000", "1011101000000000",
			"1011101000000000", "1011101000000000", "1011110000000000", "1011110000000000",
			"1011110000000000", "1011110000000000", "1011110000000000", "1011110000000000",
			"1011110000000000", "1011110000000000", "1011011010000000", "1011011010000000",
			"1011011010000000", "1011011010000000", "1011011010000000", "1011011010000000",
			"1011011010000000", "1011101000000000", "1011101000000000", "1011011000000000",
			"1011101000000000", "1011101000000000", "1011101000000000", "1011110000000000",
			"1011110000000000", "1011110000000000", "1011110000000000", "1011110000000000",
			"1011110000000000", "1011110000000000", "1011110000000000", "1011011010000000",
			"1011011010000000", "1011011010000000", "1011011010000000", "1011011010000000",
			"1011011010000000", "1011011010000000", "1011101000000000", "1011101000000000",
			"1011011000000000", "1011101000000000", "1011101000000000", "1011101000000000",
			"1011110000000000", "1011110000000000", "1011110000000000", "1011110000000000",
			"1011110000000000", "1011110000000000", "1011110000000000", "1011110000000000");

begin

	process (x)
	begin
		if (to_integer(unsigned(x) >= 6) then
			outp <= "0011110000000000";
		elsif (to_integer(unsigned(x) <= 58) then
			outp <= "1011110000000000";
		else
			outp <= tanh_lookups(to_integer(unsigned(x)));
		end if;
	end process;

end arc_hard;
