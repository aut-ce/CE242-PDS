--/*
--**********************************************************
--  Design Automation Course Homework (Spring, 2020 Semester)
--  Amirkabir University of Technology (Tehran Polytechnic)
--  Department of Computer Engineering (CE-AUT)
--  https://ce.aut.ac.ir
--  Designed TA (ali[dot]mohammadpour[at]ac[dot]ir)
--  *******************************************************
--  Student ID  : XXXXXXX
--  Student Name: -----------------
--  Student Mail: -----------------
--  *******************************************************
--  Module: ProblemSet 2, Problem 2
--  *******************************************************
--  Additional Comments:
--*/

library ieee;
use ieee.std_logic_1164.all;

entity problem_2_2 is
	port (
		a : in std_logic_vector(7 downto 0) ;
		b : in std_logic_vector(7 downto 0) ;
		c : in std_logic_vector(7 downto 0) ;
		d : in std_logic_vector(7 downto 0) ;
		mode : in std_logic ;
		y0 : out std_logic_vector(7 downto 0) ;
		y1 : out std_logic_vector(7 downto 0) ;
		y2 : out std_logic_vector(7 downto 0) ;
		y3 : out std_logic_vector(7 downto 0)) ;

end problem_2_2;

architecture problem_2_2_arc of problem_2_2 is

begin

     -- write your code here

end  problem_2_2_arc;

------------------------------------------------
------- describe new modules here --------------
------------------------------------------------
