--/*
--**********************************************************
--  Design Automation Course Homework (Spring, 2020 Semester)
--  Amirkabir University of Technology (Tehran Polytechnic)
--  Department of Computer Engineering (CE-AUT)
--  https://ce.aut.ac.ir
--  Created by TA (ali[dot]mohammadpour[at]ac[dot]ir)
--  *******************************************************
--  Student ID  : XXXXXXX
--  Student Name: -----------------
--  Student Mail: -----------------
--  *******************************************************
--  Module: ProblemSet 6, Problem 2, MAtrix Determinant
--  *******************************************************
--  Additional Comments:
--*/


entity det_matrix is
	port (
		clk : in  std_logic;
		a   : in  std_logic_vector(7 downto 0);
		b   : in  std_logic_vector(7 downto 0);
		c   : in  std_logic_vector(7 downto 0);
		d   : in  std_logic_vector(7 downto 0);
		e   : in  std_logic_vector(7 downto 0);
		f   : in  std_logic_vector(7 downto 0);
		g   : in  std_logic_vector(7 downto 0);
		h   : in  std_logic_vector(7 downto 0);
		i   : in  std_logic_vector(7 downto 0);
		det : out std_logic_vector(7 downto 0));

end det_matrix;

architecture det_matrix_arch of det_matrix is

begin

end det_matrix_arch;
