--/*
--**********************************************************
--  Design Automation Course Homework (Spring, 2020 Semester)
--  Amirkabir University of Technology (Tehran Polytechnic)
--  Department of Computer Engineering (CE-AUT)
--  https://ce.aut.ac.ir
--  Designed TA (ali[dot]mohammadpour[at]ac[dot]ir)
--  *******************************************************
--  Student ID  : XXXXXXX
--  Student ID  : XXXXXXX
--  Student Name: -----------------
--  Student Name: -----------------
--  Student Mail: -----------------
--  Student Mail: -----------------
--  *******************************************************
--  Module: PDS Project : PDS Utilities Package
--  *******************************************************
--  Additional Comments:
--*/

package pds_utils is

end package pds_utils;

package body pds_utils is

end package body pds_utils;
